LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY R_REG IS
    PORT( RST : IN  STD_LOGIC;
          CLK : IN  STD_LOGIC;
          DI  : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
          DO  : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
          RE  : IN  STD_LOGIC);
END R_REG;

ARCHITECTURE BEHAVIORAL OF R_REG IS

SIGNAL DATA : STD_LOGIC_VECTOR (15 DOWNTO 0);

BEGIN
	PROCESS(CLK, RST, RE, DATA)
	BEGIN
		IF (RST = '1') THEN
			DO <= X"0000";
			DATA <= X"0000";
		ELSIF (CLK'EVENT AND CLK = '1') THEN
			DATA <= DI;
		END IF;
		IF (RE = '1') THEN
			DO <= DATA;
		ELSE
			DO <= "ZZZZZZZZZZZZZZZZ";
		END IF;
	END PROCESS;

END BEHAVIORAL;