LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ALU IS
	GENERIC( DATA_WIDTH      : INTEGER := 15; -- DEFINING THE DATA WIDTH
		     FLAG_DATA_WIDTH : INTEGER := 3); -- DEFINING THE DATA WIDTH
	PORT( OPCODE_IN  : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		  ALU_ENABLE : IN  STD_LOGIC;
		  AIN 		 : IN  STD_LOGIC_VECTOR(DATA_WIDTH DOWNTO 0);
		  BIN        : IN  STD_LOGIC_VECTOR(DATA_WIDTH DOWNTO 0);
		  OUTP       : OUT STD_LOGIC_VECTOR(DATA_WIDTH DOWNTO 0);
		  FLAG_IN    : IN  STD_LOGIC_VECTOR(FLAG_DATA_WIDTH DOWNTO 0);
		  FLAG_OUT   : OUT STD_LOGIC_VECTOR(FLAG_DATA_WIDTH DOWNTO 0)); -- 3-V, 2-C, 1-Z, 0-S
END ALU;

ARCHITECTURE BEHAVIORAL OF ALU IS

	SIGNAL CMP_TEMP      : STD_LOGIC_VECTOR(DATA_WIDTH DOWNTO 0);
	SIGNAL YOUT 	     : STD_LOGIC_VECTOR(DATA_WIDTH DOWNTO 0);
	SIGNAL FLAG_OUT_TEMP : STD_LOGIC_VECTOR(FLAG_DATA_WIDTH DOWNTO 0);

BEGIN
	OUTP <= YOUT;
	PROCESS(AIN, BIN, OPCODE_IN, ALU_ENABLE, YOUT, CMP_TEMP, FLAG_IN, FLAG_OUT_TEMP)

		PROCEDURE FLAG_REG_CONTROL(
			AIN  : IN STD_LOGIC_VECTOR(DATA_WIDTH DOWNTO 0);
			BIN  : IN STD_LOGIC_VECTOR(DATA_WIDTH DOWNTO 0);
			YOUT : IN STD_LOGIC_VECTOR(DATA_WIDTH DOWNTO 0)) IS	
		BEGIN
			IF(YOUT = X"0000") THEN FLAG_OUT(1) <= '1';
				ELSE FLAG_OUT(1) <= '0';
			END IF;
			IF(((AIN(DATA_WIDTH) XOR BIN(DATA_WIDTH)) = '0') AND (AIN(DATA_WIDTH) = (NOT YOUT(DATA_WIDTH)))) THEN
				FLAG_OUT(3) <= '1';
			ELSE FLAG_OUT(3) <= '0';
			END IF;
			FLAG_OUT(0) <= YOUT(DATA_WIDTH);
		END PROCEDURE;
		
		PROCEDURE LOGIC_FLAG_REG_CONTROL(
			AIN  : IN STD_LOGIC_VECTOR(DATA_WIDTH DOWNTO 0);
			BIN  : IN STD_LOGIC_VECTOR(DATA_WIDTH DOWNTO 0);
			YOUT : IN STD_LOGIC_VECTOR(DATA_WIDTH DOWNTO 0)) IS	
		BEGIN
			IF(YOUT = X"0000") THEN FLAG_OUT(1) <= '1';
				ELSE FLAG_OUT(1) <= '0';
			END IF;
			FLAG_OUT(0) <= YOUT(DATA_WIDTH);
			FLAG_OUT(3) <= '0';
			FLAG_OUT(2) <= '0';
		END PROCEDURE;
		
		VARIABLE AIN_INT, BIN_INT, YOUT_INT, CARRY_TEMP_INT : INTEGER := 0;
		
	BEGIN
		CASE ALU_ENABLE IS
			WHEN '0' =>
				CASE OPCODE_IN IS
					-- NOT ENABLED
					WHEN OTHERS => NULL;
				END CASE;
			WHEN '1' =>
				AIN_INT := TO_INTEGER(UNSIGNED(AIN));
				BIN_INT := TO_INTEGER(UNSIGNED(BIN));
				CASE OPCODE_IN IS

					WHEN "0000" => -- ADD
						YOUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(AIN_INT + BIN_INT,DATA_WIDTH + 1));
						IF(AIN_INT + BIN_INT > 65535) THEN
							FLAG_OUT(2) <= '1';
						ELSE FLAG_OUT(2) <= '0';
						END IF;
						FLAG_REG_CONTROL(AIN, BIN, YOUT);

					WHEN "0001" =>	-- SUB
						IF(BIN_INT > AIN_INT) THEN YOUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(BIN_INT - AIN_INT,DATA_WIDTH + 1));
						ELSE  YOUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(AIN_INT - BIN_INT,DATA_WIDTH + 1));
						END IF;
						FLAG_OUT(2) <= '0'; --CF = 0 IF NO BORROW
						FLAG_REG_CONTROL(AIN, BIN, YOUT);

					WHEN "0010" =>	-- AND
						YOUT <= AIN AND BIN;
						LOGIC_FLAG_REG_CONTROL(AIN, BIN, YOUT);

					WHEN "0011" =>	-- OR
						YOUT <= AIN OR BIN;
						LOGIC_FLAG_REG_CONTROL(AIN, BIN, YOUT);
					
					WHEN "0100" =>	-- NOT OF BIN
						YOUT <= NOT BIN;
						
					WHEN "0101" =>	-- XOR
						YOUT <= AIN XOR BIN;
						LOGIC_FLAG_REG_CONTROL(AIN, BIN, YOUT);

					WHEN "0110" =>	-- CMP -- (BIN - AIN)
						CMP_TEMP <= STD_LOGIC_VECTOR(TO_SIGNED(BIN_INT - AIN_INT,DATA_WIDTH + 1));
						IF(BIN_INT > AIN_INT) THEN 
							FLAG_OUT(2) <= '0';
							FLAG_OUT_TEMP(2) <= '0';
						ELSE 
							FLAG_OUT(2) <= '1'; --CF = 0 IF NO BORROW
							FLAG_OUT_TEMP(2) <= '1';
						END IF;
						IF(CMP_TEMP = X"0000") THEN FLAG_OUT(1) <= '1';
						ELSE 
							FLAG_OUT(1) <= '0';
							FLAG_OUT_TEMP(1) <= '0';
						END IF;
						IF(((AIN(DATA_WIDTH) XOR BIN(DATA_WIDTH)) = '0') AND (AIN(DATA_WIDTH) = (NOT CMP_TEMP(DATA_WIDTH)))) THEN
							FLAG_OUT(3) <= '1';
							FLAG_OUT_TEMP(3) <= '1';
						ELSE 
							FLAG_OUT(3) <= '0';
							FLAG_OUT_TEMP(3) <= '0';
						END IF;
						FLAG_OUT(0) <= CMP_TEMP(DATA_WIDTH);
						FLAG_OUT_TEMP(0) <= CMP_TEMP(DATA_WIDTH);
						YOUT <= X"000" & FLAG_OUT_TEMP;


					WHEN "0111" =>	-- SHL OF BIN
						FLAG_OUT(2) <= BIN(DATA_WIDTH);
						YOUT <= STD_LOGIC_VECTOR(SHIFT_LEFT(UNSIGNED(BIN),1));
						IF((BIN(DATA_WIDTH) XOR YOUT(DATA_WIDTH)) = '1') THEN FLAG_OUT(3) <= '1';
						ELSE FLAG_OUT(3) <= '0';
						END IF;
						IF(YOUT = X"0000") THEN FLAG_OUT(1) <= '1';
						ELSE FLAG_OUT(1) <= '0';
						END IF;
						FLAG_OUT(0) <= YOUT(DATA_WIDTH);

					WHEN "1000" =>	-- SHR OF BIN
						FLAG_OUT(2) <= BIN(0);
						YOUT <= STD_LOGIC_VECTOR(SHIFT_RIGHT(UNSIGNED(BIN),1));
						IF((BIN(DATA_WIDTH) XOR YOUT(DATA_WIDTH)) = '1') THEN FLAG_OUT(3) <= '1';
						ELSE FLAG_OUT(3) <= '0';
						END IF;
						IF(YOUT = X"0000") THEN FLAG_OUT(1) <= '1';
						ELSE FLAG_OUT(1) <= '0';
						END IF;
						FLAG_OUT(0) <= YOUT(DATA_WIDTH);

					WHEN "1001" =>	-- INC OF BIN
						YOUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(BIN_INT + 1,DATA_WIDTH + 1));
						FLAG_REG_CONTROL(X"0001", BIN, YOUT);
						IF(BIN(DATA_WIDTH) = YOUT(DATA_WIDTH)) THEN FLAG_OUT(3) <= '0';
						ELSE FLAG_OUT(3) <= '1';
						END IF;

					WHEN "1010" =>	-- DEC OF BIN
						YOUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(BIN_INT - 1,DATA_WIDTH + 1));
						FLAG_REG_CONTROL(X"0001", BIN, YOUT);
						IF(BIN(DATA_WIDTH) = YOUT(DATA_WIDTH)) THEN FLAG_OUT(3) <= '0';
						ELSE FLAG_OUT(3) <= '1';
						END IF;
					
					WHEN "1011" =>	-- ROR OF BIN
					   FLAG_OUT(2) <= BIN(0);
						YOUT <= BIN(0) & BIN(DATA_WIDTH DOWNTO 1);
						IF((BIN(DATA_WIDTH) XOR YOUT(DATA_WIDTH)) = '1') THEN FLAG_OUT(3) <= '1'; -- OF = 0 IF BIN KEEPS ITS SIGN AFTER THE OPERATION
						ELSE FLAG_OUT(3) <= '0';
						END IF;
						IF(YOUT = X"0000") THEN FLAG_OUT(1) <= '1';
						ELSE FLAG_OUT(1) <= '0';
						END IF;
						FLAG_OUT(0) <= YOUT(DATA_WIDTH);
					
					WHEN "1100" =>	-- ROL OF BIN
					   FLAG_OUT(2) <= BIN(DATA_WIDTH);
						YOUT <=  BIN(DATA_WIDTH-1 DOWNTO 0) & BIN(DATA_WIDTH);
						IF((BIN(DATA_WIDTH) XOR YOUT(DATA_WIDTH)) = '1') THEN FLAG_OUT(3) <= '1'; -- OF = 0 IF BIN KEEPS ITS SIGN AFTER THE OPERATION
						ELSE FLAG_OUT(3) <= '0';
						END IF;
						IF(YOUT = X"0000") THEN FLAG_OUT(1) <= '1';
						ELSE FLAG_OUT(1) <= '0';
						END IF;
						FLAG_OUT(0) <= YOUT(DATA_WIDTH);
					
					WHEN "1101" =>	-- ADC 
						IF(FLAG_IN(2) = '1') THEN CARRY_TEMP_INT := 1;
						ELSE CARRY_TEMP_INT := 0;
						END IF;
					    YOUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(AIN_INT + BIN_INT + CARRY_TEMP_INT,DATA_WIDTH + 1));
						IF(AIN_INT + BIN_INT + CARRY_TEMP_INT > 65535) THEN
							FLAG_OUT(2) <= '1';
						ELSE FLAG_OUT(2) <= '0';
						END IF;
						FLAG_REG_CONTROL(AIN, BIN, YOUT); -- ADD WITH CARRY
						
					WHEN "1110" =>	-- SBB
						IF(BIN_INT > AIN_INT) THEN YOUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(BIN_INT - AIN_INT,DATA_WIDTH + 1));
						ELSE  YOUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(AIN_INT - BIN_INT,DATA_WIDTH + 1));
						END IF;
						FLAG_OUT(2) <= '0'; -- CF = 0 
						FLAG_REG_CONTROL(AIN, BIN, YOUT);
					
					WHEN "1111" => --MOD OF BIN
						IF (AIN_INT > 0) THEN 
							YOUT <= STD_LOGIC_VECTOR(TO_UNSIGNED(BIN_INT MOD AIN_INT,DATA_WIDTH + 1));
							FLAG_OUT(2) <= '0'; -- CF = 0, FOR MODULUS OPERATION
							FLAG_REG_CONTROL(AIN, BIN, YOUT);
						END IF;		
		
					WHEN OTHERS => NULL;
					
				END CASE;
			WHEN OTHERS => NULL;
		END CASE;
	END PROCESS;
END BEHAVIORAL;