LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY GPREG_FILE IS
    PORT( RX_W : IN    STD_LOGIC_VECTOR(13 DOWNTO 0);
          RX_R : IN    STD_LOGIC_VECTOR(13 DOWNTO 0);
          CLK  : IN    STD_LOGIC;
          RST  : IN    STD_LOGIC;
          DATA : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END GPREG_FILE;

ARCHITECTURE STRUCTURAL OF GPREG_FILE IS

  COMPONENT RW_REGISTER IS
      PORT( RST  : IN    STD_LOGIC;
            CLK  : IN    STD_LOGIC;
            DATA : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            RE   : IN    STD_LOGIC;
            WE   : IN    STD_LOGIC);
  END COMPONENT;

BEGIN

  REG0    :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(0),  RX_W(0));
  REG1    :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(1),  RX_W(1));
  REG2    :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(2),  RX_W(2));
  REG3    :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(3),  RX_W(3));
  REG4    :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(4),  RX_W(4));
  REG5    :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(5),  RX_W(5));
  REG6    :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(6),  RX_W(6));
  REG7    :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(7),  RX_W(7));
  REG8    :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(8),  RX_W(8));
  REG9    :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(9),  RX_W(9));
  REG10   :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(10), RX_W(10));
  REG11   :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(11), RX_W(11));
  REG12   :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(12), RX_W(12));
  REG13   :   RW_REGISTER     PORT MAP (RST, CLK, DATA, RX_R(13), RX_W(13));

END STRUCTURAL;