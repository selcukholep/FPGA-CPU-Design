LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BUFF IS
    PORT( PORT1	: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0); -- CPU_OUT
		  PORT2	: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0); -- CPU_IN
          RE	: IN    STD_LOGIC;
          WE	: IN    STD_LOGIC);
END BUFF;

ARCHITECTURE BEHAVIORAL OF BUFF IS
BEGIN
	PROCESS(PORT1, PORT2, RE, WE)
		BEGIN
		IF (RE = '1') THEN
			PORT2 <= PORT1;
		ELSIF(WE = '1') THEN
			PORT1 <= PORT2;
		ELSE
			PORT1 <= "ZZZZZZZZZZZZZZZZ";
			PORT2 <= "ZZZZZZZZZZZZZZZZ";
		END IF;	
	END PROCESS;
END BEHAVIORAL;