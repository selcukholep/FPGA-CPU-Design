LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FR IS
    PORT( RST : IN  STD_LOGIC;
          CLK : IN  STD_LOGIC;
          DI  : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
          DO  : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END FR;

ARCHITECTURE BEHAVIORAL OF FR IS

SIGNAL DATA : STD_LOGIC_VECTOR (3 DOWNTO 0);

BEGIN
PROCESS(CLK, RST, DATA)
BEGIN
	IF (RST = '1') THEN
		DO <= X"0";
		DATA <= X"0";
	ELSIF (CLK'EVENT AND CLK = '1') THEN
		DATA <= DI;
	END IF;
	DO <= DATA;
END PROCESS;
END BEHAVIORAL;