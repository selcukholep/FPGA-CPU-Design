LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY W_REG IS
    PORT( RST : IN  STD_LOGIC;
          CLK : IN  STD_LOGIC;
          DI  : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
          DO  : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
          WE  : IN  STD_LOGIC);
END W_REG;

ARCHITECTURE BEHAVIORAL OF W_REG IS

SIGNAL DATA : STD_LOGIC_VECTOR(15 DOWNTO 0);

BEGIN
	PROCESS(CLK, RST, WE, DI, DATA)
	BEGIN
		IF (RST = '1') THEN
			DATA <= X"0000";
			DO <= X"0000";
		ELSIF (WE = '1') THEN
			IF (CLK'EVENT AND CLK = '1') THEN
				DATA <= DI;
			END IF;
		END IF;
		DO <= DATA;
	END PROCESS;

END BEHAVIORAL;