LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY PC IS
    GENERIC( ADR_HI : STD_LOGIC_VECTOR(15 DOWNTO 0) := X"FEFF";
			 ADR_LO	: STD_LOGIC_VECTOR(15 DOWNTO 0) := X"0000");
	PORT( RST  : IN  STD_LOGIC;
          CLK  : IN  STD_LOGIC;
          WE   : IN  STD_LOGIC;
          RE   : IN  STD_LOGIC;
          UP   : IN  STD_LOGIC;
          DATA : INOUT  STD_LOGIC_VECTOR(15 DOWNTO 0));
END PC;

ARCHITECTURE BEHAVIORAL OF PC IS

SIGNAL DATA_TEMP : STD_LOGIC_VECTOR (15 DOWNTO 0);

BEGIN
	PROCESS(CLK, RST, WE, RE, UP, DATA, DATA_TEMP)
	BEGIN
		IF (RST = '1') THEN
			DATA <= ADR_LO;
			DATA_TEMP <= ADR_LO;
		ELSIF (WE = '1' OR UP = '1') THEN
			IF (CLK'EVENT AND CLK = '1') THEN
				IF (UP = '1' AND DATA_TEMP < ADR_HI) THEN
					DATA_TEMP <= STD_LOGIC_VECTOR(UNSIGNED(DATA_TEMP) + 1);
				ELSIF (DATA_TEMP = ADR_HI) THEN
					DATA_TEMP <= ADR_LO;
					DATA <= ADR_LO;
				ELSE
					DATA_TEMP <= DATA;
				END IF;
			END IF;
			DATA <= "ZZZZZZZZZZZZZZZZ";
		ELSIF (RE = '1') THEN
				DATA <= DATA_TEMP;
		ELSE
			DATA <= "ZZZZZZZZZZZZZZZZ";
		END IF;
	END PROCESS;

END BEHAVIORAL;