LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY CU IS
    PORT( RESET  : IN  STD_LOGIC;
          CLOCK  : IN  STD_LOGIC;
          IR 	   : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
          FR 	   : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
          PC_R	 : OUT STD_LOGIC;
		  		PC_U	 : OUT STD_LOGIC;
		  		PC_W	 : OUT STD_LOGIC;
		  		MAR_W	 : OUT STD_LOGIC;
		  		IR_W	 : OUT STD_LOGIC;
		  		ALU_E	 : OUT STD_LOGIC;
		  		ATR_W	 : OUT STD_LOGIC;
		  		ACC_R	 : OUT STD_LOGIC;
		  		FR_CLK : OUT STD_LOGIC;
		  		TR_W	 : OUT STD_LOGIC;
		  		TR_R	 : OUT STD_LOGIC;
		  		RX_R	 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
		  		RX_W	 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
		  		SP_R	 : OUT STD_LOGIC;
		  		SP_U	 : OUT STD_LOGIC;
		  		SP_D	 : OUT STD_LOGIC;
		  		RAM_R	 : OUT STD_LOGIC;
		  		RAM_W	 : OUT STD_LOGIC;
		  		RIO_R	 : OUT STD_LOGIC;
		  		RIO_W	 : OUT STD_LOGIC;
		  		FR_R	 : OUT STD_LOGIC;
		  		FR_W	 : OUT STD_LOGIC);
END CU;

ARCHITECTURE BEHAVIORAL OF CU IS

	COMPONENT STEPPER IS
	    PORT( CLOCK : IN  STD_LOGIC;
	          RESET : IN  STD_LOGIC := '0';
	          X     : IN  STD_LOGIC := '0';
	          Y     : IN  STD_LOGIC := '0';
	          Z     : IN  STD_LOGIC := '0';
	          W     : IN  STD_LOGIC := '0';
	          Q     : IN  STD_LOGIC := '0';
	          S     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT DECODER_4X16 IS
	    PORT( X  : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
	          Y  : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	          EN : IN  STD_LOGIC);
	END COMPONENT;
	
	SIGNAL S_RESET, X, Y, Z, W, Q : STD_LOGIC;
	SIGNAL S 					  : STD_LOGIC_VECTOR(7 DOWNTO 0); 
	SIGNAL CUD_E, SRC_E, DST_E    : STD_LOGIC;
	SIGNAL DST_BITS               : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL CUD, SRC, DST, DST2    : STD_LOGIC_VECTOR(15 DOWNTO 0);
	
	TYPE INSTRUCTION_TYPE IS (ADD_0, SUB_0, AND_0, OR_0, NOT_0, XOR_0, CMP_0, SHL_0, SHR_0, INC_0, DEC_0, ROR_0, ROL_0, ADC_0, SBB_0, MDL_0, MOV_0, XCHG_0, JMP_0, JZ_0, JNZ_0, JG_0, JLE_0, NONE_0, PUSH_0, POP_0, PUSHF_0, POPF_0, IN_0, OUT_0, NOP_0, HLT_0);
	SIGNAL INSTRUCTION : INSTRUCTION_TYPE;
	
BEGIN

	SETUP_PORTS: PROCESS(IR, RESET, CLOCK, S)
	BEGIN
		S_RESET <= RESET OR (IR(15) AND IR(14) AND IR(13) AND IR(12) AND IR(11));
		X <= (IR(7) AND IR(6) AND IR(5)) OR (IR(3) AND IR(2) AND IR(1)) OR (IR(15) AND IR(8));
		Y <= (IR(7) AND IR(6) AND IR(5) AND IR(4)) OR (IR(3) AND IR(2) AND IR(1) AND IR(0));
		Z <= (NOT IR(15)) OR (IR(15) AND IR(14) AND (NOT IR(13))) OR (IR(15) AND (NOT IR(14)) AND (NOT IR(13)) AND (NOT IR(12)) AND IR(11));
		W <= IR(15) AND IR(14) AND (NOT IR(11));
		Q <= IR(15) AND IR(8);
		
		CUD_E <= IR(15) AND (S(7) OR S(6) OR S(5));
		SRC_E <= S(7) OR S(6) OR S(5) OR (S(4) AND (NOT IR(9)));
		DST_E <= S(7) OR S(6) OR S(5) OR (S(4) AND IR(9));
	END PROCESS SETUP_PORTS;

	STEPPER_0    : STEPPER		PORT MAP(CLOCK, S_RESET, X, Y, Z, W, Q, S);
	CUD_DECODER  : DECODER_4X16	PORT MAP(IR(14 DOWNTO 11), CUD, CUD_E);
	SRC_DECODER  : DECODER_4X16	PORT MAP(IR(3 DOWNTO 0), SRC, SRC_E);
	DST_DECODER  : DECODER_4X16	PORT MAP(IR(7 DOWNTO 4), DST, DST_E);

	DST_BITS <= '0' & IR(10 DOWNTO 8);

	DST2_DECODER : DECODER_4X16	PORT MAP(DST_BITS, DST2, '1');

	PROCESS(CLOCK, RESET, S, CUD, SRC, DST, IR, FR, Z, W)
	BEGIN
		PC_U   <= S(1) OR S(3);
		PC_R   <= S(0) OR S(2);
		PC_W   <= CUD(2) OR (CUD(3) AND FR(1)) OR (CUD(4) AND (NOT FR(1))) OR (CUD(5) AND (NOT FR(2))) OR (CUD(6) AND (FR(2) OR FR(1)));
		
		MAR_W  <= S(0) OR S(2) OR S(4) OR (S(5) AND (CUD(8) OR CUD(10))) OR (S(6) AND (CUD(9) OR CUD(11)));
		IR_W   <= S(1);
		
		ALU_E  <= NOT IR(15);
		ATR_W  <= S(5) AND (NOT IR(15));
		ACC_R  <= S(7) AND (NOT IR(15));
		
		FR_CLK <= S(6) AND (NOT IR(15)) AND (NOT CLOCK);
		
		TR_W   <= S(3) OR (S(5) AND CUD(1));
		TR_R   <= (S(4) AND (NOT IR(8))) OR (SRC(14) AND ((CUD(0) AND (NOT IR(8))) OR CUD(2) OR CUD(3) OR CUD(4) OR CUD(5) OR CUD(6) OR CUD(13) OR (S(6) AND (NOT IR(15))))) OR (S(7) AND CUD(1));
		
		FOR I IN 13 DOWNTO 0 LOOP
			RX_R(I) <= (SRC(I) AND ((CUD(0) AND (NOT IR(8))) OR CUD(13) OR (S(6) AND (NOT CUD(9)) AND ( NOT CUD(10)) AND (NOT CUD(11))) OR (S(4) AND IR(8) AND (NOT IR(9))) OR (S(5) AND IR(15) AND IR(8) AND IR(9)))) OR (DST(I) AND ((S(5) AND ((NOT IR(15)) OR CUD(1))) OR (S(4) AND IR(8) AND IR(9))));
			RX_W(I) <= (DST(I) AND ((CUD(0) AND (NOT IR(8))) OR CUD(12) OR (S(7) AND DST2(7) AND (NOT IR(15)) AND (IR(14) OR (NOT IR(13)) OR (NOT IR(12)) OR IR(11))) OR (S(6) AND CUD(1)) OR (S(7) AND CUD(9)) OR (CUD(0) AND IR(8) AND (NOT IR(9))))) OR (SRC(I) AND S(7) AND CUD(1)) OR (S(7) AND (NOT IR(15)) AND DST2(I) AND (NOT DST2(7)));
		END LOOP;
		
		SP_R  <= (S(5) AND (CUD(8) OR CUD(10))) OR (S(6) AND (CUD(9) OR CUD(11)));
		SP_U  <= S(5) AND (CUD(9) OR CUD(11));
		SP_D  <= S(6) AND (CUD(8) OR CUD(10));
	
		RAM_R <= S(1) OR S(3) OR (SRC(15) AND ((CUD(0) AND (NOT IR(8))) OR CUD(13) OR (S(6) AND (NOT IR(15))))) OR (DST(15) AND (NOT IR(15)) AND S(5)) OR (S(7) AND (CUD(9) OR CUD(11))) OR (CUD(0) AND IR(8) AND (NOT IR(9)));
		RAM_W <= (DST(15) AND (CUD(0) OR CUD(12) OR (S(7) AND (NOT IR(15)) AND (IR(14) OR (NOT IR(13)) OR (NOT IR(12)) OR IR(11))))) OR (S(6) AND (CUD(8) OR CUD(10))) OR (CUD(0) AND IR(8) AND IR(9));
		
		RIO_R <= S(5) AND CUD(12);
		RIO_W <= S(5) AND CUD(13);
		
		FR_R  <= S(6) AND CUD(10);
		FR_W  <= S(7) AND CUD(11);
	
		IF ( IR(15) /= 'Z' ) THEN
			INSTRUCTION <= INSTRUCTION_TYPE'VAL(TO_INTEGER(UNSIGNED(IR(15 DOWNTO 11))));
		ELSE
			INSTRUCTION <= NONE_0;
		END IF;
	END PROCESS;

END BEHAVIORAL;