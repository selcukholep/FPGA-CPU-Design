LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY RW_REGISTER IS
    PORT( RST  : IN    STD_LOGIC;
          CLK  : IN    STD_LOGIC;
          DATA : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
          RE   : IN    STD_LOGIC;
          WE   : IN    STD_LOGIC);
END RW_REGISTER;

ARCHITECTURE BEHAVIORAL OF RW_REGISTER IS

SIGNAL DATA_TEMP : STD_LOGIC_VECTOR (15 DOWNTO 0);

BEGIN
	PROCESS(CLK, RST, RE, WE, DATA_TEMP)
	BEGIN
		IF (RST = '1') THEN
			DATA <= X"0000";
		ELSIF (WE = '1') THEN
			IF (CLK'EVENT AND CLK = '1') THEN
				DATA_TEMP <= DATA;
			END IF;
			DATA <= "ZZZZZZZZZZZZZZZZ";
		ELSIF (RE = '1') THEN
			DATA <= DATA_TEMP;
		ELSE
			DATA <= "ZZZZZZZZZZZZZZZZ";
		END IF;
	END PROCESS;

END BEHAVIORAL;