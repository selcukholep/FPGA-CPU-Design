LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY RAM IS
	GENERIC( BITS 		: INTEGER := 16 ; -- NUMBER OF BITS PER RAM WORD
			 ADDR_BITS	: INTEGER := 4 ); -- 2 ^ADDR_BITS = NUMBER OF WORDS IN RAM
	PORT( CLK  : IN    STD_LOGIC;
		  RST  : IN    STD_LOGIC;									-- RESET
		  WE   : IN    STD_LOGIC;									-- WRITE ENABLE
		  RE   : IN    STD_LOGIC;									-- READ ENABLE
		  A    : IN    STD_LOGIC_VECTOR(ADDR_BITS - 1 DOWNTO 0);	-- ADDRESS
		  DATA : INOUT STD_LOGIC_VECTOR(BITS - 1 DOWNTO 0));		-- DATA BUS
END RAM;

ARCHITECTURE BEHAVIORAL OF RAM IS

	TYPE RAM_TYPE IS ARRAY (2**ADDR_BITS - 1 DOWNTO 0 ) OF STD_LOGIC_VECTOR (BITS - 1 DOWNTO 0 );
	SIGNAL RAM : RAM_TYPE;
	SIGNAL READ_A : STD_LOGIC_VECTOR(ADDR_BITS - 1 DOWNTO 0 );

BEGIN
	PROCESS(CLK, RST, A, RE, WE, READ_A, DATA, RAM)
	BEGIN
		READ_A <= A;
		IF (RST = '1') THEN
			FOR I IN 0 TO 2**ADDR_BITS - 1 LOOP
				RAM(I) <= X"0000";
			END LOOP;
			DATA <= X"0000";
		ELSIF (WE = '1') THEN
			IF (CLK'EVENT AND CLK = '1') THEN
				RAM(CONV_INTEGER(UNSIGNED(A))) <= DATA;
			END IF;
			DATA <= "ZZZZZZZZZZZZZZZZ";
		ELSIF (RE = '1') THEN
				DATA <= RAM(CONV_INTEGER(UNSIGNED(READ_A)));
		ELSIF (RE = '0') THEN
				DATA <= "ZZZZZZZZZZZZZZZZ";
		END IF;
	END PROCESS;	

END BEHAVIORAL;