LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY IR IS
    PORT( RST : IN  STD_LOGIC;
          CLK : IN  STD_LOGIC;
          DI  : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
          DO  : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
          WE  : IN  STD_LOGIC);
END IR;

ARCHITECTURE BEHAVIORAL OF IR IS
BEGIN
	PROCESS(CLK, RST, DI, WE)
	BEGIN
		IF (RST = '1') THEN
			DO <= "ZZZZZZZZZZZZZZZZ";
		ELSIF (CLK'EVENT AND CLK = '1') THEN
			IF (WE = '1') THEN
				DO <= DI;
			END IF;
		END IF;
	END PROCESS;
END BEHAVIORAL;