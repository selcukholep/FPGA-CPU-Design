LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY CONTROLLER IS
    PORT( RESET    : IN  STD_LOGIC;
          CLOCK    : IN  STD_LOGIC;
		  TMP_DATA : INOUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		  TMP_ADR : IN	STD_LOGIC_VECTOR(15 DOWNTO 0);
		  START	   : IN  STD_LOGIC);
END CONTROLLER;

ARCHITECTURE BEHAVIORAL OF CONTROLLER IS

COMPONENT CPU IS
    PORT( RESET : IN    STD_LOGIC;
           CLOCK : IN    STD_LOGIC;
           RAM	 : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
           RAM_R : OUT   STD_LOGIC;
           RAM_W : OUT   STD_LOGIC;
		   IO	 : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		   ADR	 : OUT   STD_LOGIC_VECTOR(15 DOWNTO 0));
END COMPONENT;

COMPONENT RAM IS
	GENERIC( BITS 	   : INTEGER := 16  ;
			 ADDR_BITS : INTEGER := 16 );
	PORT( CLK  : IN    STD_LOGIC;
		  RST  : IN    STD_LOGIC;									-- RESET
		  WE   : IN    STD_LOGIC;									-- WRITE ENABLE
		  RE   : IN    STD_LOGIC;									-- READ ENABLE
		  A    : IN    STD_LOGIC_VECTOR(ADDR_BITS - 1 DOWNTO 0);	-- ADDRESS
		  DATA : INOUT STD_LOGIC_VECTOR(BITS - 1 DOWNTO 0));		-- DATA BUS
END COMPONENT;

SIGNAL CPU_RESET, CPU_RAM_R, CPU_RAM_W, RAM_W, RAM_CLOCK : STD_LOGIC;
SIGNAL CPU_RAM_ADR, IO  								 : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL RAM_ADR 											 : STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');

BEGIN

TMP_RAM_INIT : PROCESS(RESET, CLOCK, START, CPU_RAM_ADR, TMP_ADR, RAM_ADR)
	BEGIN 
		IF (START = '0') THEN
			RAM_CLOCK <= CLOCK;
		END IF;
		IF (START = '1') THEN
			RAM_ADR <= CPU_RAM_ADR;
			RAM_CLOCK <= NOT CLOCK;
		ELSIF (TMP_ADR(0) /= 'Z') THEN
			RAM_ADR <= TMP_ADR;
		ELSIF (CLOCK'EVENT AND CLOCK = '0' AND START = '0' AND RESET = '0') THEN
			RAM_ADR <= STD_LOGIC_VECTOR(UNSIGNED(RAM_ADR) + 1);
		END IF;
	END PROCESS TMP_RAM_INIT;

CPU_RESET <= NOT START;
RAM_W 	 <= CPU_RAM_W OR (NOT START);

CPU_0 : CPU PORT MAP(CPU_RESET, CLOCK, TMP_DATA, CPU_RAM_R, CPU_RAM_W, IO, CPU_RAM_ADR);
RAM_0 : RAM PORT MAP(RAM_CLOCK, RESET, RAM_W, CPU_RAM_R, RAM_ADR, TMP_DATA);

END BEHAVIORAL;
