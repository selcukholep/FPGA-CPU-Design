LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FLAG_BUFFER IS
	GENERIC( FLAG_WIDTH : INTEGER := 4 );
    PORT( PORT1	: INOUT STD_LOGIC_VECTOR(FLAG_WIDTH - 1 DOWNTO 0);
	      PORT2	: INOUT STD_LOGIC_VECTOR(FLAG_WIDTH - 1 DOWNTO 0); 
          RE	: IN    STD_LOGIC;
          WE	: IN    STD_LOGIC);
END FLAG_BUFFER;
ARCHITECTURE BEHAVIORAL OF FLAG_BUFFER IS
BEGIN
	PROCESS(PORT1, PORT2, RE, WE)
	BEGIN
		IF (RE = '1') THEN
			PORT2 <= PORT1;
		ELSIF (WE = '1') THEN
			PORT1 <= PORT2;
		ELSE
			PORT1 <= "ZZZZ";
			PORT2 <= "ZZZZ";
		END IF;
	END PROCESS;
END BEHAVIORAL;